module 
	Xor_and_gate(input a, input b, input c,  output y);
    	assign y = (a^b) & c;
endmodule
