//`timescale 1ns / 1ps
////////////////////////////////////////////////////////////////////////////////////
//// Company: 
//// Engineer: 
//// 
//// Create Date: 06/30/2025 11:38:04 AM
//// Design Name: 
//// Module Name: tb_full_adder
//// Project Name: 
//// Target Devices: 
//// Tool Versions: 
//// Description: 
//// 
//// Dependencies: 
//// 
//// Revision:
//// Revision 0.01 - File Created
//// Additional Comments:
//// 
////////////////////////////////////////////////////////////////////////////////////


//module tb_full_adder;
//    reg A, B, Cin;
//    wire Sum, Carry;

//    full_adder uut(.A(A), .B(B), .Cin(Cin), .Sum(Sum), .Carry(Carry) );

//    integer i;

//    initial begin
//    for(i = 0; i < 8; i = i+1)
//    begin
//        {A, B, Cin} = i;
//        #10;
//    end
//    $finish;
//    end        
//endmodule
