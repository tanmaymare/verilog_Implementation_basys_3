//`timescale 1ns / 1ps
////////////////////////////////////////////////////////////////////////////////////
//// Company: 
//// Engineer: 
//// 
//// Create Date: 06/24/2025 03:26:24 PM
//// Design Name: 
//// Module Name: half_adder
//// Project Name: 
//// Target Devices: 
//// Tool Versions: 
//// Description: 
//// 
//// Dependencies: 
//// 
//// Revision:
//// Revision 0.01 - File Created
//// Additional Comments:
//// 
////////////////////////////////////////////////////////////////////////////////////


//module half_adder(
//    input A,
//    input B,
//    output Sum,
//    output Carry
//);
//    assign Sum = A ^ B;
//    assign Carry = A & B;
//endmodule
